// Copyright (c) 2025 Sigma Logic

package lvds_pkg;

    typedef struct packed {
        logic p;
        logic n;
    } pair_t;

endpackage : lvds_pkg
